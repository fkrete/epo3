l
2
