l
2
mk
